module test_rx();







endmodule
